--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   02:28:00 11/22/2022
-- Design Name:   
-- Module Name:   E:/programming1/VHDL/FPU/test_sm2c.vhd
-- Project Name:  FPP
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: SM2C
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY test_sm2c IS
END test_sm2c;
 
ARCHITECTURE behavior OF test_sm2c IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT SM2C
    PORT(
         num : IN  std_logic_vector(23 downto 0);
         sign : IN  std_logic;
         numc : OUT  std_logic_vector(28 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal num : std_logic_vector(23 downto 0) := (others => '0');
   signal sign : std_logic := '0';

 	--Outputs
   signal numc : std_logic_vector(28 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
   
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: SM2C PORT MAP (
          num => num,
          sign => sign,
          numc => numc
        );
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
		
		num <= "000011110000111100101011";
		sign <= '0';
		
      wait for 100 ns;	
		
		num <= "000011110000010100100011";
		sign <= '1';		

      wait;
   end process;

END;
